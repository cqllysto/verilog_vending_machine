`timescale 1ps/1ps

module main(
    input d,n,
    output z,c
);




endmodule


